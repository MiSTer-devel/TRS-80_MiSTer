//
// HT1080Z for MiSTer IOCTL Loader Module
//
// Copyright (c) 2020 Stephen Eddy
//
// All rights reserved
//
// Redistribution and use in source and synthezised forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// * Redistributions of source code must retain the above copyright notice,
//   this list of conditions and the following disclaimer.
//
// * Redistributions in synthesized form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.
//
// * Neither the name of the author nor the names of other contributors may
//   be used to endorse or promote products derived from this software without
//   specific prior written agreement from the author.
//
// * License is granted for non-commercial use only.  A fee may not be charged
//   for redistributions as source code or in synthesized/hardware form without 
//   specific prior written agreement from the author.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
// THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
// PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.

module cmd_loader
#( parameter
        DATA = 8,                           // Data bus width
        ADDR = 16                           // Address bus width
)
(
    input wire clock, reset,                // I/O clock and async reset

    input wire      ioctl_download,         // Signal indicating an active download in progress
	input wire  [7:0]       ioctl_index,    // Menu index used to upload the file
	input wire              ioctl_wr,       // Signal be ioctl to write data (receive)
	input wire [DATA-1:0]   ioctl_dout,     // Data being sent into the loader by ioctl
	output logic            ioctl_wait,     // Signal from the laoder to hold the current output data

    output logic loader_wr,			        // Signal to write to ram
    output logic loader_download,	        // Download in progress (active high)
    output logic [ADDR-1:0] loader_addr,    // Address in ram to write data to
    output logic [DATA-1:0] loader_data,    // Data to write to ram
    output logic [ADDR-1:0] execute_addr,   // Start address for program start
    output logic execute_enable   	        // Jump to start address (out_execute_addr) - Not implemented
); 

typedef enum bit [2:0] {IDLE, GET_TYPE, GET_LEN, GET_LSB, GET_MSB, SETUP, TRANSFER, IGNORE} loader_states;
loader_states state;

always_ff @(posedge clock or posedge reset)
begin
	logic [8:0] block_len;
	logic [7:0] block_type;
	logic [15:0] block_addr;
	logic old_download;
	logic first_block;

	if (reset)
	begin
		execute_enable <= 0;
		loader_addr <= '0;
		execute_addr <= '0;
		loader_data <= '0;
		old_download <= 0;
		state <= IDLE;
		loader_download <= 0;
		ioctl_wait <= 0;
		block_addr <= '0;
	end 
	else begin

		loader_wr <= '0;
		ioctl_wait <= '0;
		execute_enable <= 0;

		case(state)
			IDLE: begin 		// No transfer occurring
				if(~old_download && ioctl_download && ioctl_index > 1) begin
					loader_download <= 1;
					state <= GET_TYPE;
				end
			end
			GET_TYPE: begin		// Start of transfer, load block type
				ioctl_wait <= 0;
				if(ioctl_wr) begin
					block_type <= ioctl_dout;
					if(ioctl_dout ==8'd0) begin	// EOF
						loader_download <= 0;
						state <= IDLE;
                    end else state <= GET_LEN;
				end
			end
			GET_LEN: begin		// Setup len or finish transfer
				if(ioctl_wr) begin
					if(block_type == 8'd1) begin
						case(ioctl_dout)
						8'd2: block_len <= 9'd256;
						8'd1: block_len <= 9'd0;
						default: block_len <= ((ioctl_dout - 2 ) & 9'd255);
						endcase
						state <= GET_LSB;
					end else if(block_type == 8'd2) begin
						block_len <= 9'd0;
						state <= GET_LSB;
					end else begin
						block_len <= ioctl_dout;
						state <= IGNORE;
					end
				end
			end
			GET_LSB: begin
				if(ioctl_wr) begin
					block_addr[7:0] <= ioctl_dout;
					state <= GET_MSB;
				end 
			end
			GET_MSB: begin
				if(ioctl_wr) begin
					block_addr[15:8] <= ioctl_dout;
					ioctl_wait <= 1;
					state <= SETUP;
				end 
			end
			SETUP: begin		
				if(block_type == 8'd1) begin	// Data block
					loader_addr <= block_addr;
					state <= TRANSFER;
				end if(block_type == 8'd2) begin	
					execute_addr <= block_addr;
					execute_enable <= 1;	// toggle execute flag
					if(block_len > 2)  begin
						state <= IGNORE; 
					end else begin
						loader_download <= 0;
						state <= IDLE; 
					end					
				end else begin	// Shoudl only ever be 1 or 2, so error state
					loader_download <= 0;
					state <= IDLE;
				end
			end
			TRANSFER: begin
				if(ioctl_wr) begin
					if(block_len > 0) begin
						loader_addr <= loader_addr + 1;
						block_len <= block_len - 1;
						loader_data <= ioctl_dout;
						loader_wr <= 1;
					end else begin	// Move to next block in chain
						state <= GET_TYPE;
						loader_wr <= 0;
					end
				end
			end
			IGNORE: begin
				if(ioctl_wr) begin
					if(block_len > 0) begin
						block_len <= block_len - 1;
					end else begin
						if(block_type == 8'd0 || block_type == 8'd2) begin
							state <= IDLE; 
							loader_download <= 0;
						end else state <= GET_TYPE;
					end
				end
			end
		endcase
        // Reset back when ioctl download ends
        if(old_download && ~ioctl_download && ioctl_index > 1) begin
            loader_download <= 0;
        end
	end
end
endmodule

